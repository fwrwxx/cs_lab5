library verilog;
use verilog.vl_types.all;
entity mux5to1_4bit_tb is
end mux5to1_4bit_tb;
